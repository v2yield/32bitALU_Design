`timescale 1ns / 1ps
module Or_32bit(
    input [31:0] a,
    input [31:0] b,
    output [31:0] s
    );

or a1 (s[0],a[0],b[0]);
or a2 (s[1],a[1],b[1]);
or a3 (s[2],a[2],b[2]);
or a4 (s[3],a[3],b[3]);
or a5 (s[4],a[4],b[4]);
or a6 (s[5],a[5],b[5]);
or a7 (s[6],a[6],b[6]);
or a8 (s[7],a[7],b[7]);
or a9 (s[8],a[8],b[8]);
or a10 (s[9],a[9],b[9]);
or a11 (s[10],a[10],b[10]);
or a12 (s[11],a[11],b[11]);
or a13 (s[12],a[12],b[12]);
or a14 (s[13],a[13],b[13]);
or a15 (s[14],a[14],b[14]);
or a16 (s[15],a[15],b[15]);
or a17 (s[16],a[16],b[16]);
or a18 (s[17],a[17],b[17]);
or a19 (s[18],a[18],b[18]);
or a20 (s[19],a[19],b[19]);
or a21 (s[20],a[20],b[20]);
or a22 (s[21],a[21],b[21]);
or a23 (s[22],a[22],b[22]);
or a24 (s[23],a[23],b[23]);
or a25 (s[24],a[24],b[24]);
or a26 (s[25],a[25],b[25]);
or a27 (s[26],a[26],b[26]);
or a28 (s[27],a[27],b[27]);
or a29 (s[28],a[28],b[28]);
or a30 (s[29],a[29],b[29]);
or a31 (s[30],a[30],b[30]);
or a32 (s[31],a[31],b[31]);

endmodule

