`timescale 1ns / 1ps
module Not_32bit(
    input [31:0] a,
    output [31:0] s
    );
    
not a1 (s[0],a[0]);
not a2 (s[1],a[1]);
not a3 (s[2],a[2]);
not a4 (s[3],a[3]);
not a5 (s[4],a[4]);
not a6 (s[5],a[5]);
not a7 (s[6],a[6]);
not a8 (s[7],a[7]);
not a9 (s[8],a[8]);
not a10 (s[9],a[9]);
not a11 (s[10],a[10]);
not a12 (s[11],a[11]);
not a13 (s[12],a[12]);
not a14 (s[13],a[13]);
not a15 (s[14],a[14]);
not a16 (s[15],a[15]);
not a17 (s[16],a[16]);
not a18 (s[17],a[17]);
not a19 (s[18],a[18]);
not a20 (s[19],a[19]);
not a21 (s[20],a[20]);
not a22 (s[21],a[21]);
not a23 (s[22],a[22]);
not a24 (s[23],a[23]);
not a25 (s[24],a[24]);
not a26 (s[25],a[25]);
not a27 (s[26],a[26]);
not a28 (s[27],a[27]);
not a29 (s[28],a[28]);
not a30 (s[29],a[29]);
not a31 (s[30],a[30]);
not a32 (s[31],a[31]);

endmodule

